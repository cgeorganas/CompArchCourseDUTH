`ifdef MODEL_TECH
	`include "../sys_defs.vh"
`endif

module fpu_flt2int(
	input	logic	[31:0]	in,
	input	logic			is_signed,
	output	logic	[34:0]	out
);



endmodule
